//`ifndef COMMON_VH
//`define COMMON_VH

`timescale 1ns/1ps

/*
-------------------------------------------------------------------------------------------------------------------
Version:
    1.5.0: 2023-05-24
           Vivado 2022.1
           Updated VERSION macro.
           RISCV cores version 1.3.2.
           Decoupled system version 2.0.2.
           Removed old video subsystem.
    
    1.5.1: 2023-06-16
           RISCV cores version 1.3.3.
           Decoupled system version 2.0.3.
           
    1.5.2: 2023-06-26
           Bootloader firmware with 100MHz system clock configuration.
           2023-06-07
           Fixed some synthesis warnings.
           2023-06-29
           Profiler for residual coding.           
    1.5.3: 2023-06-30
           Vivado 2022.2
           Fixed some Methodology critical warnings / warnings.
           2023-07-07
           Integrated HLS long tail functions.
           2023-07-13
           Integrated mtDMA for each riscv.
    1.5.4: 2023-07-14
           New DRP PLL for XMII RX   
           2023-07-18
           Updated mtDMA.
    1.5.5: 2023-08-02
           Updated from So's XMII clock.
           Updated HLS long tail functions.
           2023-08-03
           Integrated with fill_reference_samples.
           xmem interface (AXIS->xmem) for pixel_add_hls with row/column convertor.
           2023-08-04
           output pixel HLS to copy recon pixel to ddr (via cache).
           2023-08-09
           ASYNC_REG for XMII cross-clock domain register between shifted clock and non-shfited clock.
           DONT_TOUCH for HLS (intraFilter, intraPred, quant, dequant, dct, idct, getRes, pixadd).
           Fill_ref_sample HLS generated by vitis 2020.
           2023-08-10
	       Remove all DONT_TOUCH.
           2023-08-14
	       Fixed all errors reported by spyglass.
           2023-08-15
	       Fixed all warnings reported by spyglass.
           2023-08-16
           Use new riscv xmem interface with byte-write-enable.
           2023-08-22
           Macro to enable/desable XMII.
           2023-08-24
           ASYNC_OUT=0 for encodeBin/decodeBin AXI4 arbiter.
           Fixed some modelSim warnings.
           Use UI_SYSCLK from MIG instead of sysPll
           Seperate reset for m_axi_clk and system_clk
           2023-08-29
           Rollback to not using MIG output system clock.
           2023-09-05
           Rollback to use rstn to reset AXI4 256 to 512 convertor.
           Xmem with top/left pixel buffer for fill_ref_samples.
           2023-09-06
           Connect UI_RST to AXI4 256 to 512 convertor but no reset synchronizer.
           2023-09-20
           Fixed the bug of residual coding unpacker with output busy signal
           Fixed the bug of rcStream control of recon pixel.
           2023-09-21
           Added recon rc done to return queue.
           2023-09-25
           unpacker busy signal depends on tf_empty.
           2023-09-26
           Update rbsp HLS.
           Removed unused mark_debug.
           2023-09-27
           Fixed the bug of rbsp HLS integration.
           Fixed the modelSim warning about rbsp AXIS DMA.
           Riscv profilier with 32 function.
           Increase the size of FLOW_FDEC_DDR.
           2023-09-28
           Output pins for profiling functions.
           4 outpix HLS with 4 flow cache to DDR.
		   2023-11-22
		   Updated from Github.
           2023-11-29
           Cabac decoder read xmem parameter directly.
           fill_ref_sample calcluates row/buffer pointer.
           add_pixel's row-to-cow module calculate row/buffer pointer.
		   2023-12-01
		   Merged with So's K7 version
           2023-12-07
           Optimized fill_ref_sample.
           Optimized residual coding with spq without software polling done.
           Get cabac if dataflow HLS is disabled.
           2023-12-12
           Updated with So's longtail HLS.
           2023-12-14
           Each tile has its own sqp in residual coding.
           2024-01-06
           Non-blocking hls ap control interface.
           Non-blocking mtdma.
           mtdma is located before data_bus_arbiter (rollbacked on 2024-01-17).
           2024-01-09
           csr mcycle is used for cycle profiling excluded cache miss.
           2024-01-11
           fill_ref_samples write to dataflow cache directly.
		   2024-01-12
		   reduce xmem read latency.
		   2024-01-16
		   Updated with So's longtail HLS.
           Reduce decodeBin latency by 2.
           2024-01-18
           Parameter to enable longtail HLS or dataflow HLS for each core.
           For flow cache, use simple datamem instead of cache memory.
           Disable some data HLS if only decoder enabled.
           2024-01-22
           Extran return queue for CMDR dependence.
           2024-01-23
           8 outpix HLS.
           2024-01-25
           Fixed timing path of ready signal from flow cache arbiter.
           2024-01-26
           Parameter for outpix HLS number.
           2024-02-01
           Updated with Git by So.
           Added bullet riscv for testing.
    1.6.0  2024-02-05
           Testing version for bullet riscv.
           Bus interface for mutex cache.
           Bus interface for commander.
           remove BITMEM, DEBUGGER and MPU_PROTECTION.
           2024-02-15
           Added new dmaCore to replace mtDMA.
    1.6.1  2024-03-04
           Micro thread for bullet Riscv.
           Profiler for buller Riscv.
           Added macro SYSTEM_FREQUENCY.
           2024-03-07
           Fixed some synthesis warnining.
           2024-03-15
           Integrated mruCache (no mesi).
    1.6.2  2024-04-12
           Updated mseiDirectory from So.
           vsRisc5_v1_5.
           Seperate bullet riscv data and io bus.
           mcache with io mapping.
    1.6.3  2024-04-25
           bullet riscv with rollback pipeline.
           new dcache arbiter with rollback interface.
           two stages dcache arbiter is used.
    1.6.4  2024-05-02
           Optimized micro thread controller.
           Integrated mesi cache with rollback.
    1.6.5  2024-05-09
           Testing mesi cache with rollback.
           Only one AXI4 port for decoupled system.
           2024-05-14
           Remove PROF_FUNC_NUM which is useless.
           Added ENABLE_PROFILER parameter.
           12-bits AXI4 ID.
           2024-05-16
           Updated openHevc longtail HLS.
           Modified generic_cache_arbiter to match HLS cache interface.
           2024-05-17
           Updated openHevc longtail HLS (git commit id: db14cdf)
    1.6.6  2024-05-24
           New system hierarchy.
    1.6.7  2024-06-05
           Vivado 2024.1
           2024-06-06
           Fixed some warnings.
           RGMII IO port not use inout since no TSI anymore.
           Map RF write to cmdr taskqueue.
           Map jump to cmdr start.
           2024-06-13
           Update openHevc HLS.
Remark:
    For RISCV/decoupled system, please refer version description in vsRisc5_vX_X.sv, hls_dataflow_system_top_vX.sv
    and hls_longtail_system_top_vX.sv.
-------------------------------------------------------------------------------------------------------------------
*/

//Test on K7 fpga
//`define K7_FPGA_TEST

//=============================================================================
//                                  Version
//=============================================================================
`define VERSION_MAJOR    1
`define VERSION_MINOR    6
`define VERSION_PATCH    7
`define VERSION_YEAR     2024
`define VERSION_MONTH    06
`define VERSION_DAY      13

//=============================================================================
//                                Default Macro
//=============================================================================
//Default parameter in riscv_top_wrap.sv
`ifndef DEFAULT_CORE_NUM
    `define DEFAULT_CORE_NUM   4
`endif
`ifndef DEFAULT_ENABLE_HLS
    `define DEFAULT_ENABLE_HLS 1
`endif
`ifndef DEFAULT_ENABLE_PROFILER
    `define DEFAULT_ENABLE_PROFILER 1
`endif

//=============================================================================
//                                ENCODE or DECODE
//=============================================================================
`define ENABLE_DEC

//=============================================================================
//                                ASIC or FPGA
//=============================================================================
`ifdef _VIVADO_
	`define FPGA
  `ifndef K7_FPGA_TEST
	`define VU19P
  `endif
`else
	`define ASIC
`endif

//=============================================================================
//                                System Frequency
//=============================================================================
`ifdef VU19P
    `define SYSTEM_FREQUENCY     100000000
`else
    `define SYSTEM_FREQUENCY      70000000
`endif

//=============================================================================
//                                HLS
//=============================================================================
//Test to enable/disable dataflow HLS
`ifndef K7_FPGA_TEST
`define DATA_FLOW_HLS
`endif
//Test to enable/disable long tail HLS
`define LONG_TAIL_HLS

//=============================================================================
//                             OTHER PERIPHERAL
//=============================================================================
`define UART_IO_2
//`define UART_IO_3
//`define SPI_IO
//`define IR_IO
`define ENABLE_GPIO
`define NO_CLK_DIV_PAD
`define BOOTUP_SPI
`define ENABLE_I2C
`define NEW_I2C

//=============================================================================
//                                 XMII TSI
//=============================================================================
`define ENABLE_XMII                        // Enable XMII
`define FPGA_XMII                          // XMII or TSI(no used now)
`define NEW_MDIO                           // define this macro to use new clocking of MDIO data out
`define XMII_RW_BYTE_SWAP                  // define it to enable xmii read or write byte swap
//`define ENABLE_XMII_DRP_PLL
//=============================================================================
//                                 Include Files
//=============================================================================
//Define Bus mapping
`include "busDefine.vh"

//=============================================================================
//                               MARCO for SOFTWARE RESET
//=============================================================================
//`define SOFT_RESET                       // define it to enable Riscv reset via csr instruction

//=============================================================================
//                               MARCO for WATCHDOG
//=============================================================================
//`define WATCHDOG                         // define it to enable Riscv watchdog via csr instruction

//=============================================================================
//                               MARCO for AXILITE_DRP
//=============================================================================
//`define AXILITE_DRP                      // define it to enable AXILITE DRP MMCM
//`define TEST_BRAM2AXILITE_MASTER         // define it only for SIMULATION of the riscv_to_axilite_master module with axilite bram device
                                           // default please remove this macro define for normal operation

//=============================================================================
//                             MACRO FOR MQSTAT
//=============================================================================
`define MQSTAT


//=============================================================================
//                               MARCO for VESA SUBSYSTEM
//=============================================================================

//Enable vesa_subsystem
`define ENABLE_VESA


//=============================================================================
//                               MARCO for XMEM
//=============================================================================
`define ENABLE_OPENHEVC


//=============================================================================
//                            AXI4_DATA_WIDTH_CONV MARCO used by So
//=============================================================================
`define AXI_DWIDTH_CONV_SYNC_FIFO_NAME axi_dwidth_conv_sync_fifo
