// Decode Bin Interface
always_comb begin
    decBin_get_c = '{default:'0};
    decBin_ctx_c = '{default:'0};
    decBin_sel_c = '{default:'0};

${statement}
end
